----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:16:55 04/11/2010 
-- Design Name: 
-- Module Name:    fakecogram - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity fakecogram is
	port (
		clka: IN std_logic;
		dina: IN std_logic_VECTOR(31 downto 0);
		addra: IN std_logic_VECTOR(8 downto 0);
		wea: IN std_logic_VECTOR(0 downto 0);
		douta: OUT std_logic_VECTOR(31 downto 0);
		clkb: IN std_logic;
		dinb: IN std_logic_VECTOR(31 downto 0);
		addrb: IN std_logic_VECTOR(8 downto 0);
		web: IN std_logic_VECTOR(0 downto 0);
		doutb: OUT std_logic_VECTOR(31 downto 0)
	);
end fakecogram;

architecture Behavioral of fakecogram is
	signal stuff	: std_logic_vector(16383 downto 0)	:= 
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"00000000000000000000000000000000" &
"11111111111111111111111111111111" &	-- -1
"01011100011111000000000000000111" &	--jmp #7
"10100111101111000001000000001000" &	--neg 8, 8		--should give -2
"01101111111111000001000000001000" &	--xor 8, #8		--should give 2
"01100011111111000001000000001111" &	--and 8, #0xF	--should give A
"01101011111111000001000010101010" &	--or 8, #0xAA	--should give AA
"10000111111111000001000000000010" &	--sub 8, #2		--should give 0
"10000011111111000001000000000001" &	--add 8, #1		--should give 2
"10101011101111000001000000001000";		--abs 8, 8		--should give 1
	signal aa	: integer;
	signal ab	: integer;
begin
	aa <= to_integer(unsigned(addra));
	ab <= to_integer(unsigned(addrb));

	process(clka)
	begin
		if rising_edge(clka) then
			if wea(0)='1' then
				stuff(aa*32+31 downto aa*32) <= dina;
			else
				douta <= stuff(aa*32+31 downto aa*32);
			end if;
		end if;
	end process;
	
	process(clkb)
	begin
		if rising_edge(clkb) then
			doutb <= stuff(ab*32+31 downto ab*32);
		end if;
	end process;
end Behavioral;

